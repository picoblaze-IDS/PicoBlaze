----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:39:10 12/02/2010 
-- Design Name: 
-- Module Name:    CPU_and_Table - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity CPU_and_Table is
    PORT(

         match_strobe : OUT  std_logic;
         out_port : OUT  std_logic_vector(7 downto 0);
         interrupt : IN  std_logic;
         interrupt_ack : OUT  std_logic;
         reset : IN  std_logic;
         clk : IN  std_logic
        );
end CPU_and_Table;

architecture Behavioral of CPU_and_Table is

    -- Component Declaration for the processor and its program store
 
    COMPONENT embedded_kcpsm3
    PORT(
         port_id : OUT  std_logic_vector(7 downto 0);
         write_strobe : OUT  std_logic;
         read_strobe : OUT  std_logic;
         out_port : OUT  std_logic_vector(7 downto 0);
         in_port : IN  std_logic_vector(7 downto 0);
         interrupt : IN  std_logic;
         interrupt_ack : OUT  std_logic;
         reset : IN  std_logic;
         clk : IN  std_logic
        );
    END COMPONENT;

--
-- declaration of the data table
--

component dataTable is
    Generic(
	     -- port address, for picoblaze
		  -- Note: set this to an EVEN value.
        portnumber : std_logic_vector(7 downto 0);
		  
       INIT_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"

    ); 
    Port (
        CLK : in  STD_LOGIC;
        RST : in std_logic;
        RD : in  STD_LOGIC;
        WR : in  STD_LOGIC;
        PORT_ID : in  STD_LOGIC_VECTOR (7 downto 0);
        DATA_IN : in std_logic_vector (7 downto 0);
        DATA_OUT : out  STD_LOGIC_VECTOR (7 downto 0) );
end component;

signal port_id : std_logic_vector(7 downto 0);
signal write_strobeI : std_logic;
signal out_portI : std_logic_vector(7 downto 0);
signal read_strobe : std_logic;
signal in_port : std_logic_vector(7 downto 0);

signal src0 : std_logic_vector(7 downto 0);
signal src1 : std_logic_vector(7 downto 0);

constant MATCHPORTNUMBER : std_logic_vector(7 downto 0) := "00001000";
signal SEL : std_logic;

begin

	-- Instantiate the processor and its program store
   uut: embedded_kcpsm3 PORT MAP (
        port_id => port_id,
        write_strobe => write_strobeI,
        read_strobe => read_strobe,
        out_port => out_portI,
        in_port => in_port,
        interrupt => interrupt,
        interrupt_ack => interrupt_ack,
        reset => reset,
        clk => clk );
		  
    -- when we output to MATCHPORTNUMBER, then the data will be on out_port and
	 -- the match_strobe signal will go to logic 1.
    out_port <= out_portI;
    SEL <= '1' when PORT_ID(7 downto 0)=MATCHPORTNUMBER(7 downto 0) else '0';	 
    match_strobe <= write_strobeI AND SEL;
	
    -- match data	table
    dt: dataTable
	 generic map
	 (
	     portnumber => "00000100",
		  
        -- each INIT line has 32 bytes, which are arranged in order *right to left*
        -- hence the following line has the values 0 to 31 in order of increasing value
        -- INIT_00 => "1F1E1D1C1B1A191817161514131211100F0E0D0C0B0A09080706050403020100",
		  
INIT_00 => X"2400620100000000000000025C01730108016D018400650118002F0100000000",
INIT_01 => X"00000000000000033C006E010000000000000003300069010000000000000003",
INIT_02 => X"5C01000360006801000000001800000354007301000000000000000348002F01",
INIT_03 => X"1501A8C01501A8C0FFFF0000FFFFFFFF00000000060000040000000301000000",
INIT_04 => X"00000000000000039C0074010000000000000003900078010000000016001600",
INIT_05 => X"08010003C0006F010000000000000003B4006D010000000000000003A8002001",
INIT_06 => X"E40074010000000020010003D8006E010000000014010003CC00750100000000",
INIT_07 => X"0001A8C0FFFF0000FF01A8C00001A8C00600000438010003020000002C010003",
INIT_08 => X"0000000320017501000000000000000314016F01000000006F006F00FF01A8C0",
INIT_09 => X"0000000303000000000000033801740100000000000000032C016E0100000000",
INIT_0A => X"000000006F006F00FF01A8C00001A8C0FFFF0000FFFFFFFF0000000006000004",
INIT_0B => X"0000000380016501000000000000000374016301000000000000000368017501",
INIT_0C => X"A4016501000000000000000398016D0100000000840000038C01200100000000",
INIT_0D => X"000000005C010003BC0120010000000084000003B00173010000000008010003",
INIT_0E => X"00000003E00175010000000000000003D4016F010000000000000003C8016201",
INIT_0F => X"040273010000000000000003F80165010000000000000003EC016C0100000000",
INIT_10 => X"080706051E000A000403020104030201060000045C0100030400000084000003",
INIT_11 => X"0000000000000000000000000000000000000000000000004500450008070605"


	 )
	 port map
	 (
        CLK => clk,
        RST => reset,
        RD => read_strobe,
        WR => write_strobeI,
        PORT_ID => port_id,
        DATA_IN => out_portI,
        DATA_OUT => src0
    );
	 
	 -- network data table
	 nw: dataTable
	 generic map
	 (
	     portnumber => "00000110",
		          
        -- each INIT line has 32 bytes, which are arranged in order *right to left*
        -- hence the following line has the values 0 to 31 in order of increasing value
        -- "1F1E1D1C1B1A191817161514131211100F0E0D0C0B0A09080706050403020100"
INIT_00 => X"060504030201000006720040A96B420000450008006C3DF72400F9ACB73B1F00",
INIT_01 => X"1600E4574F040A08010100005D72FE0018803C5CCF87D18E330D450014000807",
INIT_02 => X"686571776A65207177656A207177656A71776A68656A686A7177686A7177AAA0",
INIT_03 => X"656A206B71772065686A77716B2065687177206B65776871206B656871776B20",
INIT_04 => X"71776B6820656A6B77716865206A6B777168206A656B777168206A656B717768",
INIT_05 => X"6B777120686B77712068656A6B77712068656B77716820656A6B71776820656A",
INIT_06 => X"6820656A6B77716820656A6B71776820656A6B777168206A656B77712068656A",
INIT_07 => X"6A6B77716820656A6B77716820656A6B77716820656A6B77716820656A6B7771",
INIT_08 => X"77656A71776A68656A686A7177686A717765206B77716820656A6B7771682065",
INIT_09 => X"2065687177206B65776871206B656871776B20686571776A65207177656A2071",
INIT_0A => X"6A6B777168206A656B777168206A656B717768656A206B71772065686A77716B",
INIT_0B => X"77712068656B77716820656A6B71776820656A71776B6820656A6B7771686520",
INIT_0C => X"776820656A6B777168206A656B77712068656A6B777120686B77712068656A6B",
INIT_0D => X"656A6B77716820656A6B77716820656A6B77716820656A6B77716820656A6B71",
INIT_0E => X"686A717765206B77716820656A6B77716820656A6B77716820656A6B77716820",
INIT_0F => X"656871776B20686571776A65207177656A207177656A71776A68656A686A7177",
INIT_10 => X"6A656B717768656A206B71772065686A77716B2065687177206B65776871206B",
INIT_11 => X"71776820656A71776B6820656A6B77716865206A6B777168206A656B77716820",
INIT_12 => X"77712068656A6B777120686B77712068656A6B77712068656B77716820656A6B",
INIT_13 => X"20656A6B77716820656A6B77716820656A6B71776820656A6B777168206A656B",
INIT_14 => X"6B77716820656A6B77716820656A6B77716820656A6B77716820656A6B777168",
INIT_15 => X"7177656A207177656A71776A68656A686A7177686A717765206B77716820656A",
INIT_16 => X"65686A77716B2065687177206B65776871206B656871776B20686571776A6520",
INIT_17 => X"6B77716865206A6B777168206A656B777168206A656B717768656A206B717720",
INIT_18 => X"712068656A6B77712068656B77716820656A6B71776820656A71776B6820656A",
INIT_19 => X"6820656A6B71776820656A6B777168206A656B77712068656A6B777120686B77",
INIT_1A => X"6A6B77716820656A6B77716820656A6B77716820656A6B77716820656A6B7771",
INIT_1B => X"656A686A7177686A717765206B77716820656A6B77716820656A6B7771682065",
INIT_1C => X"65776871206B656871776B20686571776A65207177656A207177656A71776A68",
INIT_1D => X"656B777168206A656B717768656A206B71772065686A77716B2065687177206B",
INIT_1E => X"716820656A6B71776820656A71776B6820656A6B77716865206A6B777168206A",
INIT_1F => X"7168206A656B77712068656A6B777120686B77712068656A6B77712068656B77",
INIT_20 => X"656A6B77716820656A6B77716820656A6B77716820656A6B71776820656A6B77",
INIT_21 => X"00000000000000000073656C756F622073656D206563757320656A6B77716820"
	 )
	 port map
	 (
        CLK => clk,
        RST => reset,
        RD => read_strobe,
        WR => write_strobeI,
        PORT_ID => port_id,
        DATA_IN => out_portI,
        DATA_OUT => src1
    );
	 
	 in_port <= src0 when port_id(2 downto 1) = "10" else
	            src1 when port_id(2 downto 1) = "11" else
					"00000000";
					
end Behavioral;

